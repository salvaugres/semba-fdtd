* dual rc ladder
R1 in 0 10
I1 0 in dc 0
.tran 50u 200u
.save v(in)
.end